** sch_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/top_level_1st_order.sch
**.subckt top_level_1st_order
x1 net2 GND net3 BJT2 BJTs
x2 VDD net1 BJT2 net2 GND CTAT
x3 VDD net1 BJT2 V GND net3 PTAT
V1 VDD GND 5
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.control
dc temp -40 125 0.1
plot v(V)
*plot v(V4,PTAT)
*let CTAT1 = v(CTAT)*i(CTAT)
*plot v(CTAT1)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  BJTs.sym # of pins=4
** sym_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/BJTs.sym
** sch_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/BJTs.sch
.subckt BJTs  BJT VSS BJT1 BJT2
*.iopin VSS
*.iopin BJT
*.iopin BJT1
*.iopin BJT2
XQ10 VSS VSS BJT sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ11 VSS VSS BJT sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ13 VSS VSS BJT sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ14 VSS VSS BJT sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ15 VSS VSS BJT sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ12 VSS VSS BJT1 sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ9 VSS VSS BJT2 sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends


* expanding   symbol:  CTAT.sym # of pins=5
** sym_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/CTAT.sym
** sch_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/CTAT.sch
.subckt CTAT  VDD PTAT V1 BJT VSS
*.iopin VDD
*.iopin PTAT
*.iopin V1
*.iopin BJT
*.iopin VSS
XM22 PTAT net3 net4 VSS sky130_fd_pr__nfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM23 net3 net3 V1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM24 net1 PTAT VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM25 net3 net4 net1 VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=30 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM26 net2 PTAT VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM29 PTAT V1 net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=30 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 BJT net4 VSS sky130_fd_pr__res_high_po_0p35 L=8 mult=1 m=1
XR2 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=8 mult=1 m=1
XR3 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=8 mult=1 m=1
.ends


* expanding   symbol:  PTAT.sym # of pins=6
** sym_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/PTAT.sym
** sch_path: /home/shahid/Desktop/EDA/test_BGR/xschem_BGR/PTAT.sch
.subckt PTAT  VDD PTAT V1 V VSS BJT1
*.iopin VDD
*.iopin PTAT
*.iopin V1
*.iopin BJT1
*.iopin V
*.iopin VSS
XM27 net1 PTAT VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM28 V V1 net1 VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=30 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR2 net2 V VSS sky130_fd_pr__res_high_po_0p35 L=44.43 mult=1 m=1
XR1 BJT1 net2 VSS sky130_fd_pr__res_high_po_0p35 L=44.43 mult=1 m=1
XR3 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=44.43 mult=1 m=1
XR4 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=44.43 mult=1 m=1
.ends

.GLOBAL GND
.end
