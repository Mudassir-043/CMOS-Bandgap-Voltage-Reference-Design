** sch_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/BGR_2ndc.sch
**.subckt BGR_2ndc Vfinal VNL V_first IBIAS VSS VDD
*.opin Vfinal
*.iopin VNL
*.iopin V_first
*.iopin IBIAS
*.iopin VSS
*.iopin VDD
XR3 Vfinal net1 VSS sky130_fd_pr__res_high_po_0p35 L=3.2 mult=1 m=1
XR4 net1 net2 VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR5 net2 net3 VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR12 net3 net4 VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR13 net4 net5 VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR14 net5 VNL VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR1 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR2 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
XR6 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=3.2 mult=1 m=1
XR7 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=3.2 mult=1 m=1
x1 VDD VSS V_first net1 Vfinal IBIAS Opamp_Jaffar_withBlocks
**.ends

* expanding   symbol:  Opamp_Jaffar_withBlocks.sym # of pins=6
** sym_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/Opamp_Jaffar_withBlocks.sym
** sch_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/Opamp_Jaffar_withBlocks.sch
.subckt Opamp_Jaffar_withBlocks  VDD VSS VP VN VO IBIAS
*.iopin VDD
*.iopin VSS
*.iopin VP
*.iopin VN
*.iopin VO
*.iopin IBIAS
x1 VSS VO IBIAS net1 Current_mirror_jaffar
x2 VDD VSS VP VN net1 VO Diff_Opamp_jaffar
XC2 VDD VSS sky130_fd_pr__cap_mim_m3_1 W=30 L=10 MF=1 m=1
XC3 VDD VSS sky130_fd_pr__cap_mim_m3_1 W=30 L=10 MF=1 m=1
.ends


* expanding   symbol:  Current_mirror_jaffar.sym # of pins=4
** sym_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/Current_mirror_jaffar.sym
** sch_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/Current_mirror_jaffar.sch
.subckt Current_mirror_jaffar  VSS VO IBIAS SO
*.iopin VSS
*.iopin VO
*.iopin IBIAS
*.iopin SO
XM2 SO IBIAS net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=50 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 VO IBIAS net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=100 nf=20 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 IBIAS IBIAS net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=50 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net2 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net3 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=100 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  Diff_Opamp_jaffar.sym # of pins=6
** sym_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/Diff_Opamp_jaffar.sym
** sch_path: /home/shahid/Desktop/EDA/test/xschem_BGR_Top/Diff_Opamp_jaffar.sch
.subckt Diff_Opamp_jaffar  VDD VSS VP VN SO VO
*.iopin VDD
*.iopin VSS
*.iopin VP
*.iopin VN
*.iopin SO
*.iopin VO
XM30 net2 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM32 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM31 net1 VN SO VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=50 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 VP SO VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=50 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 net3 VO sky130_fd_pr__cap_mim_m3_1 W=24 L=24 MF=1 m=1
XM6 VO net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=100 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 net3 net2 VSS sky130_fd_pr__res_high_po_0p35 L=8 mult=1 m=1
.ends

.end
