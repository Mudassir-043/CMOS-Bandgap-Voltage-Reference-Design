** sch_path: /home/shahid/Desktop/EDA/test/xschem BGR/BGR_2nd_partb_Mubashir.sch
**.subckt BGR_2nd_partb_Mubashir VDD VSS V2 V4 VNL
*.iopin VDD
*.iopin VSS
*.iopin V2
*.iopin V4
*.iopin VNL
XM9 net3 V4 net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=5 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net1 V2 net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 VNL net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM58 net2 VDD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=5 W=20 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR11 net3 VNL VSS sky130_fd_pr__res_high_po_0p35 L=47 mult=1 m=1
XR1 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=47 mult=1 m=1
XR2 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 L=47 mult=1 m=1
**.ends
.end
